`define SYNTHESIS
`define sfuzz_rand_reg rand reg
